module LCD (
    input i_rst,
    input i_clk,   
    
    output [7:0] o_LCD_DATA,
    output       o_LCD_EN,
    output       o_LCD_RS,
    output       o_LCD_RW,
    output       o_LCD_ON,
    output       o_LCD_BLON
);



endmodule